module spart_tb();

