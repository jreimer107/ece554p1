module spart_tb();

reg [6:0] HEX0, HEX1, HEX2, HEX3, HEX4, HEX5;
